module numpad (
	input clk;
	output [3:0]reg out
);

//bla bla bla

endmodule
