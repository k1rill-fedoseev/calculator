module display (
	input clock,
	output [7:0] ctrl,
	output [7:0] led
);

//  ###0###
// #       #
// #       #
// 5       1
// #       #
// #       #
//  ###6###
// #       #
// #       #
// 4       2
// #       # ###
// #       # #7#
//  ###3###  ###

//        76543210
//
// 0 - 8'b00111111
// 1 - 8'b00000110
// 2 - 8'b01011011
// 3 - 8'b01001111
// 4 - 8'b01100110
// 5 - 8'b01101101
// 6 - 8'b01111101
// 7 - 8'b00000111
// 8 - 8'b01111111
// 9 - 8'b01101111
// . - 8'b10000000

reg [13:0] counter = 0;

always  @(posedge clock)
begin: a1
	
end

endmodule
