module numpad (
	input clk,
	output [3:0] rows,
	input [3:0] columns,
	output [4:0] value
);

//bla bla bla

endmodule