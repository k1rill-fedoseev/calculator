module display (
input clk;
output [7:0]ctrl;
output [7:0]leds
);



endmodule
