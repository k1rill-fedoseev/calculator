module numpad (
    input clock,
    input [3:0] rows,
    output [3:0] columns,
    output [4:0] value
);

endmodule
